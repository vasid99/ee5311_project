*** SPICE deck for cell wavtest{sch} from library project_kansu3
*** Created on Sat Jan 09, 2021 18:52:17
*** Last revised on Sat Jan 09, 2021 18:53:51
*** Written on Sat Jan 09, 2021 18:53:55 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 0.1, MIN_CAPAC 0.01FF

.global gnd

*** TOP LEVEL CELL: wavtest{sch}

* Spice Code nodes in cell cell 'wavtest{sch}'
V1 A gnd wavfile="/home/vasid/.git/courses/dic_proj/spice_scripts/fa_characterize/fa_char_inputs0.wav"
.tran 0 1n
.END
