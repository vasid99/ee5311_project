*** SPICE deck for cell sta_char_and{sch} from library project_kansu3
*** Created on Sun Jan 10, 2021 14:20:35
*** Last revised on Sun Jan 10, 2021 14:22:36
*** Written on Mon Jan 11, 2021 02:45:21 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 0.1, MIN_CAPAC 0.01FF

* cell 'and1x{sch}' is described in this file:
.include /home/vasid/.git/courses/dic_proj/SPI_files/and1x.spi

* cell 'fa_c3x_s2x{sch}' is described in this file:
.include /home/vasid/.git/courses/dic_proj/SPI_files/fa_c3x_s2x.spi

*** TOP LEVEL CELL: sta_char_and{sch}
Xand1x@0 A_in B_in gnd vdd Y_out and1x
Xfa_c3x_s@0 fa_c3x_s@0_A fa_c3x_s@0_B Y_out fa_c3x_s@0_Co_bar gnd fa_c3x_s@0_S_bar vdd fa_c3x_s2x

* Spice Code nodes in cell cell 'sta_char_and{sch}'
.include "/home/vasid/.git/courses/dic_proj/spice_scripts/and_characterize/script1.txt"
.END
