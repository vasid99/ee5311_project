*** SPICE deck for cell csm_non_pipelined{sch} from library project_kansu3
*** Created on Tue Dec 22, 2020 17:35:14
*** Last revised on Sat Jan 09, 2021 10:33:41
*** Written on Sat Jan 09, 2021 10:33:42 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 0.1, MIN_CAPAC 0.01FF

*** SUBCIRCUIT project_kansu3__and1x FROM CELL and1x{sch}
.SUBCKT project_kansu3__and1x A B Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 net@13 A net@50 gnd nmos_HP L=0.022U W=0.088U
Mnmos@2 Y net@13 gnd gnd nmos_HP L=0.022U W=0.044U
Mnmos@3 net@50 B gnd gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 vdd A net@13 vdd pmos_HP L=0.022U W=0.088U
Mpmos@1 vdd B net@13 vdd pmos_HP L=0.022U W=0.088U
Mpmos@3 vdd net@13 Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project_kansu3__and1x

*** SUBCIRCUIT project_kansu3__fa_c3x_s2x FROM CELL fa_c3x_s2x{sch}
.SUBCKT project_kansu3__fa_c3x_s2x A B Ci Co_bar S_bar
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@33 B net@40 gnd nmos_HP L=0.022U W=0.132U
Mnmos@1 S_bar Ci net@33 gnd nmos_HP L=0.022U W=0.132U
Mnmos@2 net@40 A gnd gnd nmos_HP L=0.022U W=0.132U
Mnmos@3 net@21 A gnd gnd nmos_HP L=0.022U W=0.176U
Mnmos@4 net@21 B gnd gnd nmos_HP L=0.022U W=0.176U
Mnmos@5 S_bar Co_bar net@21 gnd nmos_HP L=0.022U W=0.176U
Mnmos@6 net@21 Ci gnd gnd nmos_HP L=0.022U W=0.176U
Mnmos@7 Co_bar Ci net@73 gnd nmos_HP L=0.022U W=0.264U
Mnmos@8 net@73 A gnd gnd nmos_HP L=0.022U W=0.264U
Mnmos@9 net@73 B gnd gnd nmos_HP L=0.022U W=0.264U
Mnmos@10 net@67 A gnd gnd nmos_HP L=0.022U W=0.088U
Mnmos@11 Co_bar B net@67 gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 net@20 Ci S_bar vdd pmos_HP L=0.022U W=0.264U
Mpmos@1 net@1 B net@20 vdd pmos_HP L=0.022U W=0.264U
Mpmos@2 vdd A net@1 vdd pmos_HP L=0.022U W=0.264U
Mpmos@3 net@25 Co_bar S_bar vdd pmos_HP L=0.022U W=0.352U
Mpmos@4 vdd A net@25 vdd pmos_HP L=0.022U W=0.352U
Mpmos@5 vdd B net@25 vdd pmos_HP L=0.022U W=0.352U
Mpmos@6 vdd Ci net@25 vdd pmos_HP L=0.022U W=0.352U
Mpmos@7 net@49 Ci Co_bar vdd pmos_HP L=0.022U W=0.528U
Mpmos@8 vdd A net@49 vdd pmos_HP L=0.022U W=0.528U
Mpmos@9 vdd B net@49 vdd pmos_HP L=0.022U W=0.528U
Mpmos@10 vdd A net@62 vdd pmos_HP L=0.022U W=0.176U
Mpmos@11 net@62 B Co_bar vdd pmos_HP L=0.022U W=0.176U
.ENDS project_kansu3__fa_c3x_s2x

*** SUBCIRCUIT project_kansu3__inv1x FROM CELL inv1x{sch}
.SUBCKT project_kansu3__inv1x A Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y A gnd gnd nmos_HP L=0.022U W=0.044U
Mpmos@0 vdd A Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project_kansu3__inv1x

*** SUBCIRCUIT project_kansu3__nand1x FROM CELL nand1x{sch}
.SUBCKT project_kansu3__nand1x A B Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@2 Y B net@3 gnd nmos_HP L=0.022U W=0.088U
Mnmos@4 net@3 A gnd gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 vdd B Y vdd pmos_HP L=0.022U W=0.088U
Mpmos@2 vdd A Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project_kansu3__nand1x

.global gnd vdd

*** TOP LEVEL CELL: csm_non_pipelined{sch}
Xand1x@0 x0 y0 z0 project_kansu3__and1x
Xand1x@7 x7 y0 x7y0 project_kansu3__and1x
Xand1x@15 x7 y1 x7y1 project_kansu3__and1x
Xand1x@16 x0 y2 x0y2 project_kansu3__and1x
Xand1x@17 x1 y2 x1y2 project_kansu3__and1x
Xand1x@18 x2 y2 x2y2 project_kansu3__and1x
Xand1x@19 x3 y2 x3y2 project_kansu3__and1x
Xand1x@20 x4 y2 x4y2 project_kansu3__and1x
Xand1x@21 x5 y2 x5y2 project_kansu3__and1x
Xand1x@22 x6 y2 x6y2 project_kansu3__and1x
Xand1x@31 x7 y3 x7y3 project_kansu3__and1x
Xand1x@32 x0 y4 x0y4 project_kansu3__and1x
Xand1x@33 x1 y4 x1y4 project_kansu3__and1x
Xand1x@34 x2 y4 x2y4 project_kansu3__and1x
Xand1x@35 x3 y4 x3y4 project_kansu3__and1x
Xand1x@36 x4 y4 x4y4 project_kansu3__and1x
Xand1x@37 x5 y4 x5y4 project_kansu3__and1x
Xand1x@38 x6 y4 x6y4 project_kansu3__and1x
Xand1x@47 x7 y5 x7y5 project_kansu3__and1x
Xand1x@48 x0 y6 x0y6 project_kansu3__and1x
Xand1x@49 x1 y6 x1y6 project_kansu3__and1x
Xand1x@50 x2 y6 x2y6 project_kansu3__and1x
Xand1x@51 x3 y6 x3y6 project_kansu3__and1x
Xand1x@52 x4 y6 x4y6 project_kansu3__and1x
Xand1x@53 x5 y6 x5y6 project_kansu3__and1x
Xand1x@54 x6 y6 x6y6 project_kansu3__and1x
Xand1x@56 x0 y7 x0y7 project_kansu3__and1x
Xand1x@57 x1 y7 x1y7 project_kansu3__and1x
Xand1x@58 x2 y7 x2y7 project_kansu3__and1x
Xand1x@59 x3 y7 x3y7 project_kansu3__and1x
Xand1x@60 x4 y7 x4y7 project_kansu3__and1x
Xand1x@61 x5 y7 x5y7 project_kansu3__and1x
Xand1x@62 x6 y7 x6y7 project_kansu3__and1x
Xfa_c3x_s2x@0 vdd INVx0y1 INVx1y0 FA_Co_bar_0_0 z1 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@1 vdd INVx1y1 INVx2y0 FA_Co_bar_0_1 FA_S_bar_0_1 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@2 vdd INVx2y1 INVx3y0 FA_Co_bar_0_2 FA_S_bar_0_2 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@3 vdd INVx3y1 INVx4y0 FA_Co_bar_0_3 FA_S_bar_0_3 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@4 vdd INVx4y1 INVx5y0 FA_Co_bar_0_4 FA_S_bar_0_4 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@5 vdd INVx5y1 INVx6y0 FA_Co_bar_0_5 FA_S_bar_0_5 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@6 vdd INVx6y1 x7y0 FA_Co_bar_0_6 FA_S_bar_0_6 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@7 vdd x7y1 gnd FA_Co_bar_0_7 FA_S_bar_0_7 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@8 FA_Co_bar_0_0 x0y2 FA_S_bar_0_1 FA_Co_bar_1_0 FA_S_bar_1_0 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@9 FA_Co_bar_0_1 x1y2 FA_S_bar_0_2 FA_Co_bar_1_1 FA_S_bar_1_1 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@10 FA_Co_bar_0_2 x2y2 FA_S_bar_0_3 FA_Co_bar_1_2 FA_S_bar_1_2 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@11 FA_Co_bar_0_3 x3y2 FA_S_bar_0_4 FA_Co_bar_1_3 FA_S_bar_1_3 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@12 FA_Co_bar_0_4 x4y2 FA_S_bar_0_5 FA_Co_bar_1_4 FA_S_bar_1_4 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@13 FA_Co_bar_0_5 x5y2 FA_S_bar_0_6 FA_Co_bar_1_5 FA_S_bar_1_5 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@14 FA_Co_bar_0_6 x6y2 FA_S_bar_0_7 FA_Co_bar_1_6 FA_S_bar_1_6 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@15 FA_Co_bar_0_7 INVx7y2 gnd FA_Co_bar_1_7 FA_S_bar_1_7 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@16 FA_Co_bar_1_0 INVx0y3 FA_S_bar_1_1 FA_Co_bar_2_0 z3 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@17 FA_Co_bar_1_1 INVx1y3 FA_S_bar_1_2 FA_Co_bar_2_1 FA_S_bar_2_1 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@18 FA_Co_bar_1_2 INVx2y3 FA_S_bar_1_3 FA_Co_bar_2_2 FA_S_bar_2_2 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@19 FA_Co_bar_1_3 INVx3y3 FA_S_bar_1_4 FA_Co_bar_2_3 FA_S_bar_2_3 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@20 FA_Co_bar_1_4 INVx4y3 FA_S_bar_1_5 FA_Co_bar_2_4 FA_S_bar_2_4 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@21 FA_Co_bar_1_5 INVx5y3 FA_S_bar_1_6 FA_Co_bar_2_5 FA_S_bar_2_5 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@22 FA_Co_bar_1_6 INVx6y3 FA_S_bar_1_7 FA_Co_bar_2_6 FA_S_bar_2_6 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@23 FA_Co_bar_1_7 x7y3 vdd FA_Co_bar_2_7 FA_S_bar_2_7 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@24 FA_Co_bar_2_0 x0y4 FA_S_bar_2_1 FA_Co_bar_3_0 FA_S_bar_3_0 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@25 FA_Co_bar_2_1 x1y4 FA_S_bar_2_2 FA_Co_bar_3_1 FA_S_bar_3_1 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@26 FA_Co_bar_2_2 x2y4 FA_S_bar_2_3 FA_Co_bar_3_2 FA_S_bar_3_2 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@27 FA_Co_bar_2_3 x3y4 FA_S_bar_2_4 FA_Co_bar_3_3 FA_S_bar_3_3 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@28 FA_Co_bar_2_4 x4y4 FA_S_bar_2_5 FA_Co_bar_3_4 FA_S_bar_3_4 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@29 FA_Co_bar_2_5 x5y4 FA_S_bar_2_6 FA_Co_bar_3_5 FA_S_bar_3_5 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@30 FA_Co_bar_2_6 x6y4 FA_S_bar_2_7 FA_Co_bar_3_6 FA_S_bar_3_6 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@31 FA_Co_bar_2_7 INVx7y4 gnd FA_Co_bar_3_7 FA_S_bar_3_7 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@32 FA_Co_bar_3_0 INVx0y5 FA_S_bar_3_1 FA_Co_bar_4_0 z5 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@33 FA_Co_bar_3_1 INVx1y5 FA_S_bar_3_2 FA_Co_bar_4_1 FA_S_bar_4_1 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@34 FA_Co_bar_3_2 INVx2y5 FA_S_bar_3_3 FA_Co_bar_4_2 FA_S_bar_4_2 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@35 FA_Co_bar_3_3 INVx3y5 FA_S_bar_3_4 FA_Co_bar_4_3 FA_S_bar_4_3 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@36 FA_Co_bar_3_4 INVx4y5 FA_S_bar_3_5 FA_Co_bar_4_4 FA_S_bar_4_4 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@37 FA_Co_bar_3_5 INVx5y5 FA_S_bar_3_6 FA_Co_bar_4_5 FA_S_bar_4_5 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@38 FA_Co_bar_3_6 INVx6y5 FA_S_bar_3_7 FA_Co_bar_4_6 FA_S_bar_4_6 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@39 FA_Co_bar_3_7 x7y5 vdd FA_Co_bar_4_7 FA_S_bar_4_7 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@40 FA_Co_bar_4_0 x0y6 FA_S_bar_4_1 FA_Co_bar_5_0 FA_S_bar_5_0 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@41 FA_Co_bar_4_1 x1y6 FA_S_bar_4_2 FA_Co_bar_5_1 FA_S_bar_5_1 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@42 FA_Co_bar_4_2 x2y6 FA_S_bar_4_3 FA_Co_bar_5_2 FA_S_bar_5_2 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@43 FA_Co_bar_4_3 x3y6 FA_S_bar_4_4 FA_Co_bar_5_3 FA_S_bar_5_3 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@44 FA_Co_bar_4_4 x4y6 FA_S_bar_4_5 FA_Co_bar_5_4 FA_S_bar_5_4 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@45 FA_Co_bar_4_5 x5y6 FA_S_bar_4_6 FA_Co_bar_5_5 FA_S_bar_5_5 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@46 FA_Co_bar_4_6 x6y6 FA_S_bar_4_7 FA_Co_bar_5_6 FA_S_bar_5_6 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@47 FA_Co_bar_4_7 INVx7y6 gnd FA_Co_bar_5_7 FA_S_bar_5_7 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@48 FA_Co_bar_5_0 x0y7 FA_S_bar_5_1 FA_Co_bar_6_0 z7 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@49 FA_Co_bar_5_1 x1y7 FA_S_bar_5_2 FA_Co_bar_6_1 FA_S_bar_6_1 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@50 FA_Co_bar_5_2 x2y7 FA_S_bar_5_3 FA_Co_bar_6_2 FA_S_bar_6_2 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@51 FA_Co_bar_5_3 x3y7 FA_S_bar_5_4 FA_Co_bar_6_3 FA_S_bar_6_3 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@52 FA_Co_bar_5_4 x4y7 FA_S_bar_5_5 FA_Co_bar_6_4 FA_S_bar_6_4 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@53 FA_Co_bar_5_5 x5y7 FA_S_bar_5_6 FA_Co_bar_6_5 FA_S_bar_6_5 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@54 FA_Co_bar_5_6 x6y7 FA_S_bar_5_7 FA_Co_bar_6_6 FA_S_bar_6_6 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@55 FA_Co_bar_5_7 INVx7y7 vdd FA_Co_bar_6_7 FA_S_bar_6_7 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@56 FA_Co_bar_6_0 gnd FA_S_bar_6_1 FA_Co_bar_7_0 FA_S_bar_7_0 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@57 net@2026 FA_Co_bar_7_0 net@2028 FA_Co_bar_7_1 z9 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@58 FA_Co_bar_6_2 FA_Co_bar_7_1 FA_S_bar_6_3 FA_Co_bar_7_2 FA_S_bar_7_2 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@59 net@2031 FA_Co_bar_7_2 net@2033 FA_Co_bar_7_3 z11 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@60 FA_Co_bar_6_4 FA_Co_bar_7_3 FA_S_bar_6_5 FA_Co_bar_7_4 FA_S_bar_7_4 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@61 net@2036 FA_Co_bar_7_4 net@2037 FA_Co_bar_7_5 z13 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@62 FA_Co_bar_6_6 FA_Co_bar_7_5 FA_S_bar_6_7 FA_Co_bar_7_6 FA_S_bar_7_6 project_kansu3__fa_c3x_s2x
Xfa_c3x_s2x@63 net@2040 FA_Co_bar_7_6 gnd Cdrop z15 project_kansu3__fa_c3x_s2x
Xinv@0 FA_Co_bar_6_1 net@2026 project_kansu3__inv1x
Xinv@1 FA_S_bar_6_2 net@2028 project_kansu3__inv1x
Xinv@2 FA_Co_bar_6_3 net@2031 project_kansu3__inv1x
Xinv@3 FA_S_bar_6_4 net@2033 project_kansu3__inv1x
Xinv@4 FA_Co_bar_6_5 net@2036 project_kansu3__inv1x
Xinv@5 FA_S_bar_6_6 net@2037 project_kansu3__inv1x
Xinv@6 FA_Co_bar_6_7 net@2040 project_kansu3__inv1x
Xinv@7 FA_S_bar_1_0 z2 project_kansu3__inv1x
Xinv@8 FA_S_bar_3_0 z4 project_kansu3__inv1x
Xinv@9 FA_S_bar_5_0 z6 project_kansu3__inv1x
Xinv@10 FA_S_bar_7_0 z8 project_kansu3__inv1x
Xinv@11 FA_S_bar_7_2 z10 project_kansu3__inv1x
Xinv@12 FA_S_bar_7_4 z12 project_kansu3__inv1x
Xinv@13 FA_S_bar_7_6 z14 project_kansu3__inv1x
Xnand1x@1 x1 y0 INVx1y0 project_kansu3__nand1x
Xnand1x@2 x2 y0 INVx2y0 project_kansu3__nand1x
Xnand1x@3 x3 y0 INVx3y0 project_kansu3__nand1x
Xnand1x@4 x4 y0 INVx4y0 project_kansu3__nand1x
Xnand1x@5 x5 y0 INVx5y0 project_kansu3__nand1x
Xnand1x@6 x6 y0 INVx6y0 project_kansu3__nand1x
Xnand1x@8 x0 y1 INVx0y1 project_kansu3__nand1x
Xnand1x@9 x1 y1 INVx1y1 project_kansu3__nand1x
Xnand1x@10 x2 y1 INVx2y1 project_kansu3__nand1x
Xnand1x@11 x3 y1 INVx3y1 project_kansu3__nand1x
Xnand1x@12 x4 y1 INVx4y1 project_kansu3__nand1x
Xnand1x@13 x5 y1 INVx5y1 project_kansu3__nand1x
Xnand1x@14 x6 y1 INVx6y1 project_kansu3__nand1x
Xnand1x@23 x7 y2 INVx7y2 project_kansu3__nand1x
Xnand1x@24 x0 y3 INVx0y3 project_kansu3__nand1x
Xnand1x@25 x1 y3 INVx1y3 project_kansu3__nand1x
Xnand1x@26 x2 y3 INVx2y3 project_kansu3__nand1x
Xnand1x@27 x3 y3 INVx3y3 project_kansu3__nand1x
Xnand1x@28 x4 y3 INVx4y3 project_kansu3__nand1x
Xnand1x@29 x5 y3 INVx5y3 project_kansu3__nand1x
Xnand1x@30 x6 y3 INVx6y3 project_kansu3__nand1x
Xnand1x@39 x7 y4 INVx7y4 project_kansu3__nand1x
Xnand1x@40 x0 y5 INVx0y5 project_kansu3__nand1x
Xnand1x@41 x1 y5 INVx1y5 project_kansu3__nand1x
Xnand1x@42 x2 y5 INVx2y5 project_kansu3__nand1x
Xnand1x@43 x3 y5 INVx3y5 project_kansu3__nand1x
Xnand1x@44 x4 y5 INVx4y5 project_kansu3__nand1x
Xnand1x@45 x5 y5 INVx5y5 project_kansu3__nand1x
Xnand1x@46 x6 y5 INVx6y5 project_kansu3__nand1x
Xnand1x@55 x7 y6 INVx7y6 project_kansu3__nand1x
Xnand1x@63 x7 y7 INVx7y7 project_kansu3__nand1x

* Spice Code nodes in cell cell 'csm_non_pipelined{sch}'
.include "/home/vasid/.git/courses/dic_proj/spice_scripts/pathDelayCalc/script2.txt"
.END
