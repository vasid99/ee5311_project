*** SPICE deck for cell sta_char_fa_critpath{sch} from library project_kansu3
*** Created on Sat Jan 09, 2021 18:52:17
*** Last revised on Mon Jan 11, 2021 02:41:07
*** Written on Mon Jan 11, 2021 02:41:51 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 0.1, MIN_CAPAC 0.01FF

* cell 'fa_c3x_s2x{sch}' is described in this file:
.include /home/vasid/.git/courses/dic_proj/SPI_files/fa_c3x_s2x.spi

*** TOP LEVEL CELL: sta_char_fa_critpath{sch}
XCo_bar_load Co_bar_out Co_bar_load_B Co_bar_load_Ci Co_bar_load_Co_bar gnd Co_bar_load_S_bar vdd fa_c3x_s2x
XS_bar_load S_bar_load_A S_bar_load_B S_bar_out S_bar_load_Co_bar gnd S_bar_load_S_bar vdd fa_c3x_s2x
Xdut A_in B_in Ci_in Co_bar_out gnd S_bar_out vdd fa_c3x_s2x

* Spice Code nodes in cell cell 'sta_char_fa_critpath{sch}'
.include "/home/vasid/.git/courses/dic_proj/spice_scripts/fa_characterize/script1.txt"
.END
