*** SPICE deck for cell sta_char_fa_vmerge2{sch} from library project_kansu3
*** Created on Sat Jan 09, 2021 18:52:17
*** Last revised on Sun Jan 10, 2021 21:47:43
*** Written on Mon Jan 11, 2021 02:52:42 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 0.1, MIN_CAPAC 0.01FF

* cell 'fa_c3x_s2x{sch}' is described in this file:
.include /home/vasid/.git/courses/dic_proj/SPI_files/fa_c3x_s2x.spi

* cell 'inv1x{sch}' is described in this file:
.include /home/vasid/.git/courses/dic_proj/SPI_files/inv1x.spi

*** TOP LEVEL CELL: sta_char_fa_vmerge2{sch}
Xdut A_in B_in Ci_in Co_bar_out gnd S_bar_out vdd fa_c3x_s2x
Xdut_1 dut_1_A Co_bar_out dut_1_Ci dut_1_Co_bar gnd dut_1_S_bar vdd fa_c3x_s2x
Xinv1x@0 S_bar_out gnd vdd inv1x@0_Y inv1x

* Spice Code nodes in cell cell 'sta_char_fa_vmerge2{sch}'
.include "/home/vasid/.git/courses/dic_proj/spice_scripts/vmerge_characterize/script1.txt"
.END
