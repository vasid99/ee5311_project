*** SPICE deck for cell sta_char_ff_x7{sch} from library project_kansu3
*** Created on Sun Jan 10, 2021 23:17:46
*** Last revised on Sun Jan 10, 2021 23:24:41
*** Written on Sun Jan 10, 2021 23:26:25 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 0.1, MIN_CAPAC 0.01FF

*** SUBCIRCUIT project_kansu3__and1x FROM CELL and1x{sch}
.SUBCKT project_kansu3__and1x A B Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 net@13 A net@50 gnd nmos_HP L=0.022U W=0.088U
Mnmos@2 Y net@13 gnd gnd nmos_HP L=0.022U W=0.044U
Mnmos@3 net@50 B gnd gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 vdd A net@13 vdd pmos_HP L=0.022U W=0.088U
Mpmos@1 vdd B net@13 vdd pmos_HP L=0.022U W=0.088U
Mpmos@3 vdd net@13 Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project_kansu3__and1x

*** SUBCIRCUIT project_kansu3__nand1x FROM CELL nand1x{sch}
.SUBCKT project_kansu3__nand1x A B Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@2 Y B net@3 gnd nmos_HP L=0.022U W=0.088U
Mnmos@4 net@3 A gnd gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 vdd B Y vdd pmos_HP L=0.022U W=0.088U
Mpmos@2 vdd A Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project_kansu3__nand1x

*** SUBCIRCUIT project_kansu3__inv1x FROM CELL inv1x{sch}
.SUBCKT project_kansu3__inv1x A Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y A gnd gnd nmos_HP L=0.022U W=0.044U
Mpmos@0 vdd A Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project_kansu3__inv1x

*** SUBCIRCUIT project_kansu3__Tristate FROM CELL Tristate{sch}
.SUBCKT project_kansu3__Tristate clk1 D Q
** GLOBAL gnd
** GLOBAL vdd
Mnmos@2 net@9 D gnd gnd nmos_HP L=0.022U W=0.088U
Mnmos@3 Q clk1 net@9 gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 vdd D net@8 vdd pmos_HP L=0.022U W=0.176U
Mpmos@1 net@8 clk_bar Q vdd pmos_HP L=0.022U W=0.176U
Xinv@0 clk1 clk_bar project_kansu3__inv1x
.ENDS project_kansu3__Tristate

*** SUBCIRCUIT project_kansu3__staticFF FROM CELL staticFF{sch}
.SUBCKT project_kansu3__staticFF clk1 D Y
** GLOBAL gnd
** GLOBAL vdd
XTristate@2 clk1 D net@1 project_kansu3__Tristate
XTristate@3 clk_bar net@6 net@1 project_kansu3__Tristate
XTristate@4 clk_bar net@6 net@5 project_kansu3__Tristate
XTristate@5 clk1 net@49 net@5 project_kansu3__Tristate
Xinv@1 net@1 net@6 project_kansu3__inv1x
Xinv@2 net@5 Y project_kansu3__inv1x
Xinv@3 clk1 clk_bar project_kansu3__inv1x
Xinv@4 net@5 net@49 project_kansu3__inv1x
.ENDS project_kansu3__staticFF

.global gnd vdd

*** TOP LEVEL CELL: sta_char_ff_x7{sch}
Xand1x@0 net@11 vdd x7y0 project_kansu3__and1x
Xand1x@1 net@11 vdd x7y1 project_kansu3__and1x
Xand1x@2 net@11 vdd x7y3 project_kansu3__and1x
Xand1x@3 net@11 vdd x7y5 project_kansu3__and1x
Xnand1x@0 net@11 vdd INVx7y2 project_kansu3__nand1x
Xnand1x@1 net@11 vdd INVx7y4 project_kansu3__nand1x
Xnand1x@2 net@11 vdd INVx7y6 project_kansu3__nand1x
Xnand1x@3 net@11 vdd INVx7y7 project_kansu3__nand1x
XstaticFF@0 clk1 D net@11 project_kansu3__staticFF

* Spice Code nodes in cell cell 'sta_char_ff_x7{sch}'
.include "/home/vasid/.git/courses/dic_proj/spice_scripts/ff_x7_characterize/script1.txt"
.END
