*** SPICE deck for cell sta_char_fa_vmerge1{sch} from library project_kansu3
*** Created on Sat Jan 09, 2021 18:52:17
*** Last revised on Sun Jan 10, 2021 21:47:34
*** Written on Sun Jan 10, 2021 22:01:04 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 0.1, MIN_CAPAC 0.01FF

*** SUBCIRCUIT project_kansu3__fa_c3x_s2x FROM CELL fa_c3x_s2x{sch}
.SUBCKT project_kansu3__fa_c3x_s2x A B Ci Co_bar S_bar
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@33 B net@40 gnd nmos_HP L=0.022U W=0.132U
Mnmos@1 S_bar Ci net@33 gnd nmos_HP L=0.022U W=0.132U
Mnmos@2 net@40 A gnd gnd nmos_HP L=0.022U W=0.132U
Mnmos@3 net@21 A gnd gnd nmos_HP L=0.022U W=0.176U
Mnmos@4 net@21 B gnd gnd nmos_HP L=0.022U W=0.176U
Mnmos@5 S_bar Co_bar net@21 gnd nmos_HP L=0.022U W=0.176U
Mnmos@6 net@21 Ci gnd gnd nmos_HP L=0.022U W=0.176U
Mnmos@7 Co_bar Ci net@73 gnd nmos_HP L=0.022U W=0.264U
Mnmos@8 net@73 A gnd gnd nmos_HP L=0.022U W=0.264U
Mnmos@9 net@73 B gnd gnd nmos_HP L=0.022U W=0.264U
Mnmos@10 net@67 A gnd gnd nmos_HP L=0.022U W=0.088U
Mnmos@11 Co_bar B net@67 gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 net@20 Ci S_bar vdd pmos_HP L=0.022U W=0.264U
Mpmos@1 net@1 B net@20 vdd pmos_HP L=0.022U W=0.264U
Mpmos@2 vdd A net@1 vdd pmos_HP L=0.022U W=0.264U
Mpmos@3 net@25 Co_bar S_bar vdd pmos_HP L=0.022U W=0.352U
Mpmos@4 vdd A net@25 vdd pmos_HP L=0.022U W=0.352U
Mpmos@5 vdd B net@25 vdd pmos_HP L=0.022U W=0.352U
Mpmos@6 vdd Ci net@25 vdd pmos_HP L=0.022U W=0.352U
Mpmos@7 net@49 Ci Co_bar vdd pmos_HP L=0.022U W=0.528U
Mpmos@8 vdd A net@49 vdd pmos_HP L=0.022U W=0.528U
Mpmos@9 vdd B net@49 vdd pmos_HP L=0.022U W=0.528U
Mpmos@10 vdd A net@62 vdd pmos_HP L=0.022U W=0.176U
Mpmos@11 net@62 B Co_bar vdd pmos_HP L=0.022U W=0.176U
.ENDS project_kansu3__fa_c3x_s2x

*** SUBCIRCUIT project_kansu3__inv1x FROM CELL inv1x{sch}
.SUBCKT project_kansu3__inv1x A Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Y A gnd gnd nmos_HP L=0.022U W=0.044U
Mpmos@0 vdd A Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project_kansu3__inv1x

*** SUBCIRCUIT project_kansu3__Tristate FROM CELL Tristate{sch}
.SUBCKT project_kansu3__Tristate clk1 D Q
** GLOBAL gnd
** GLOBAL vdd
Mnmos@2 net@9 D gnd gnd nmos_HP L=0.022U W=0.088U
Mnmos@3 Q clk1 net@9 gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 vdd D net@8 vdd pmos_HP L=0.022U W=0.176U
Mpmos@1 net@8 clk_bar Q vdd pmos_HP L=0.022U W=0.176U
Xinv@0 clk1 clk_bar project_kansu3__inv1x
.ENDS project_kansu3__Tristate

*** SUBCIRCUIT project_kansu3__staticFF FROM CELL staticFF{sch}
.SUBCKT project_kansu3__staticFF clk1 D Y
** GLOBAL gnd
** GLOBAL vdd
XTristate@2 clk1 D net@1 project_kansu3__Tristate
XTristate@3 clk_bar net@6 net@1 project_kansu3__Tristate
XTristate@4 clk_bar net@6 net@5 project_kansu3__Tristate
XTristate@5 clk1 net@49 net@5 project_kansu3__Tristate
Xinv@1 net@1 net@6 project_kansu3__inv1x
Xinv@2 net@5 Y project_kansu3__inv1x
Xinv@3 clk1 clk_bar project_kansu3__inv1x
Xinv@4 net@5 net@49 project_kansu3__inv1x
.ENDS project_kansu3__staticFF

.global gnd vdd

*** TOP LEVEL CELL: sta_char_fa_vmerge1{sch}
Xdut A_in B_in Ci_in Co_bar_out S_bar_out project_kansu3__fa_c3x_s2x
Xdut_1 dut_1_A Co_bar_out dut_1_Ci dut_1_Co_bar dut_1_S_bar project_kansu3__fa_c3x_s2x
XstaticFF@0 vdd S_bar_out staticFF@0_Y project_kansu3__staticFF

* Spice Code nodes in cell cell 'sta_char_fa_vmerge1{sch}'
.include "/home/vasid/.git/courses/dic_proj/spice_scripts/vmerge_characterize/script1.txt"
.END
