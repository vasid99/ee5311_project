*** SPICE deck for cell sta_char_ff_x7{sch} from library project
*** Created on Sun Jan 10, 2021 23:17:46
*** Last revised on Tue Jan 12, 2021 20:44:14
*** Written on Tue Jan 12, 2021 20:44:26 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 0.1, MIN_CAPAC 0.01FF

*** SUBCIRCUIT project__and1x FROM CELL and1x{sch}
.SUBCKT project__and1x A B gnd vdd Y
Mnmos@1 net@13 A net@50 gnd nmos_HP L=0.022U W=0.088U
Mnmos@2 Y net@13 gnd gnd nmos_HP L=0.022U W=0.044U
Mnmos@3 net@50 B gnd gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 vdd A net@13 vdd pmos_HP L=0.022U W=0.088U
Mpmos@1 vdd B net@13 vdd pmos_HP L=0.022U W=0.088U
Mpmos@3 vdd net@13 Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project__and1x

*** SUBCIRCUIT project__nand1x FROM CELL nand1x{sch}
.SUBCKT project__nand1x A B gnd vdd Y
Mnmos@2 Y B net@3 gnd nmos_HP L=0.022U W=0.088U
Mnmos@4 net@3 A gnd gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 vdd B Y vdd pmos_HP L=0.022U W=0.088U
Mpmos@2 vdd A Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project__nand1x

*** SUBCIRCUIT project__inv1x FROM CELL inv1x{sch}
.SUBCKT project__inv1x A gnd vdd Y
Mnmos@0 Y A gnd gnd nmos_HP L=0.022U W=0.044U
Mpmos@0 vdd A Y vdd pmos_HP L=0.022U W=0.088U
.ENDS project__inv1x

*** SUBCIRCUIT project__Tristate FROM CELL Tristate{sch}
.SUBCKT project__Tristate clk1 D gnd Q vdd
Mnmos@2 net@9 D gnd gnd nmos_HP L=0.022U W=0.088U
Mnmos@3 Q clk1 net@9 gnd nmos_HP L=0.022U W=0.088U
Mpmos@0 vdd D net@8 vdd pmos_HP L=0.022U W=0.176U
Mpmos@1 net@8 clk_bar Q vdd pmos_HP L=0.022U W=0.176U
Xinv@0 clk1 gnd vdd clk_bar project__inv1x
.ENDS project__Tristate

*** SUBCIRCUIT project__staticFF FROM CELL staticFF{sch}
.SUBCKT project__staticFF clk1 D gnd vdd Y
XTristate@2 clk1 D gnd net@1 vdd project__Tristate
XTristate@3 clk_bar net@6 gnd net@1 vdd project__Tristate
XTristate@4 clk_bar net@6 gnd net@5 vdd project__Tristate
XTristate@5 clk1 net@49 gnd net@5 vdd project__Tristate
Xinv@1 net@1 gnd vdd net@6 project__inv1x
Xinv@2 net@5 gnd vdd Y project__inv1x
Xinv@3 clk1 gnd vdd clk_bar project__inv1x
Xinv@4 net@5 gnd vdd net@49 project__inv1x
.ENDS project__staticFF

*** TOP LEVEL CELL: sta_char_ff_x7{sch}
Xand1x@0 Yout vdd gnd vdd x7y0 project__and1x
Xand1x@1 Yout vdd gnd vdd x7y1 project__and1x
Xand1x@2 Yout vdd gnd vdd x7y3 project__and1x
Xand1x@3 Yout vdd gnd vdd x7y5 project__and1x
Xnand1x@0 Yout vdd gnd vdd INVx7y2 project__nand1x
Xnand1x@1 Yout vdd gnd vdd INVx7y4 project__nand1x
Xnand1x@2 Yout vdd gnd vdd INVx7y6 project__nand1x
Xnand1x@3 Yout vdd gnd vdd INVx7y7 project__nand1x
XstaticFF@0 clk1 D gnd vdd Yout project__staticFF

* Spice Code nodes in cell cell 'sta_char_ff_x7{sch}'
.include "../spice_scripts/char_ff_x7.txt"
.END
